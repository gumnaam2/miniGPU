library ieee;
use ieee.std_logic_1164.all;
--
--entity mux is
--	port (x0, x1: in std_logic;
--			control: in std_logic;
--			selected: out std_logic);
--end mux;
--
--architecture muxarch of mux is
--begin
--	selected <= (x0 and not control) or (x1 and control);
--end muxarch;
